library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- usado nas flags
entity reg01bit is
    port(
        clk,wr_en,reset: in std_logic;
        data_in: in std_logic;
        data_out: out std_logic
    );
end entity;


architecture a_reg01bit of reg01bit is  
signal registro: std_logic;
begin

process(clk,wr_en,reset)
begin
    if reset = '1' then
        registro <= '0';
    elsif wr_en = '1' then
        if rising_edge(clk) then
            registro <= data_in;
        end if;
    end if;
end process;

data_out <= registro;

end architecture;