library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port (
        clk      : in std_logic;
        endereco : in unsigned(6 downto 0);
        dado     : out unsigned(17 downto 0)
    );
end entity;

architecture a_rom of rom is

    type mem is array (0 to 127) of unsigned(17 downto 0);
    constant conteudo_rom : mem := (
        
        -- --- Inicialização 
        0  => B"00000001_00_000_01_001", -- LD R0, 1
        1  => B"01101111_00_001_01_001", -- LD R1, 111
        2  => B"00100001_00_010_01_001", -- LD R2, 33
        3  => B"00000001_00_011_01_001", -- LD R3, 1
        
        -- Label Loop_Inicialização
        4  => B"000000000_000_0_00_010", -- MOV AccA, R0
        5  => B"000000000_001_0_11_001", -- SW [R1], AccA
        6  => B"000000000_000_0_00_010", -- MOV AccA, R0
        7  => B"000000000_011_0_00_011", -- ADD AccA, R3
        8  => B"000000000_000_0_01_010", -- MOV R0, AccA
        9  => B"000000000_001_0_00_010", -- MOV AccA, R1
        10 => B"000000000_011_0_00_011", -- ADD AccA, R3
        11 => B"000000000_001_0_01_010", -- MOV R1, AccA
        12 => B"000000000_000_0_00_010", -- MOV AccA, R0
        13 => B"0_1110111_0_010_0_10_101", -- CNJE R2, AccA, -9 

        -- Crivo 2 
        14 => B"01110010_00_001_01_001", -- LD R1, 114
        15 => B"00000010_00_011_01_001", -- LD R3, 2
        16 => B"00000000_00_100_01_001", -- LD R4, 0
        17 => B"01001000_00_010_01_001", -- LD R2, 72
        18 => B"000000000_010_0_00_010", -- MOV AccA, R2
        19 => B"000000000_010_0_00_011", -- ADD AccA, R2
        20 => B"000000000_010_0_01_010", -- MOV R2, AccA

        -- Label Loop_Crivo_2
        21 => B"000000000_100_0_00_010", -- MOV AccA, R4
        22 => B"000000000_001_0_11_001", -- SW [R1], AccA
        23 => B"000000000_001_0_00_010", -- MOV AccA, R1
        24 => B"000000000_011_0_00_011", -- ADD AccA, R3
        25 => B"000000000_001_0_01_010", -- MOV R1, AccA
        26 => B"0_1111011_0_010_0_10_101", -- CNJE R2, AccA, -5

        -- Crivo 3 
        27 => B"01110100_00_001_01_001", -- LD R1, 116
        28 => B"00000011_00_011_01_001", -- LD R3, 3
        29 => B"01000111_00_010_01_001", -- LD R2, 71
        30 => B"000000000_010_0_00_010", -- MOV AccA, R2
        31 => B"01001000_00_010_01_001", -- LD R2, 72
        32 => B"000000000_010_0_00_011", -- ADD AccA, R2
        33 => B"000000000_010_0_01_010", -- MOV R2, AccA
        
        -- Label Loop_Crivo_3
        34 => B"000000000_100_0_00_010", -- MOV AccA, R4
        35 => B"000000000_001_0_11_001", -- SW [R1], AccA
        36 => B"000000000_001_0_00_010", -- MOV AccA, R1
        37 => B"000000000_011_0_00_011", -- ADD AccA, R3
        38 => B"000000000_001_0_01_010", -- MOV R1, AccA
        39 => B"0_1111011_0_010_0_10_101", -- CNJE R2, AccA, -5

        -- Crivo 5
        40 => B"01111000_00_001_01_001", -- LD R1, 120
        41 => B"00000101_00_011_01_001", -- LD R3, 5
        42 => B"01001000_00_010_01_001", -- LD R2, 72
        43 => B"000000000_010_0_00_010", -- MOV AccA, R2
        44 => B"01001001_00_010_01_001", -- LD R2, 73
        45 => B"000000000_010_0_00_011", -- ADD AccA, R2
        46 => B"000000000_010_0_01_010", -- MOV R2, AccA
        
        -- Label Loop_Crivo_5
        47 => B"000000000_100_0_00_010", -- MOV AccA, R4
        48 => B"000000000_001_0_11_001", -- SW [R1], AccA
        49 => B"000000000_001_0_00_010", -- MOV AccA, R1
        50 => B"000000000_011_0_00_011", -- ADD AccA, R3
        51 => B"000000000_001_0_01_010", -- MOV R1, AccA
        52 => B"0_1111011_0_010_0_10_101", -- CNJE R2, AccA, -5

        -- Prepara para OUTPUT
        53 => B"01110000_00_001_01_001", -- LD R1, 112
        54 => B"00000001_00_011_01_001", -- LD R3, 1
        55 => B"01000111_00_010_01_001", -- LD R2, 71
        56 => B"000000000_010_0_00_010", -- MOV AccA, R2
        57 => B"01001000_00_010_01_001", -- LD R2, 72
        58 => B"000000000_010_0_00_011", -- ADD AccA, R2
        59 => B"000000000_010_0_01_010", -- MOV R2, AccA
        60 => B"00000000_00_100_01_001", -- LD R4, 0        

        -- Label Loop_Print_R5 
        61 => B"0000000_00_001_1_10_001", -- LW AccB, [R1]
        
        -- Se AccB != 0 (É Primo), Pula 2 linhas 
        62 => B"0_0000010_1_100_1_10_101", -- CNJE R4, AccB, +2
        
        -- Pula para 65 (Não colo 0 no R5)
        63 => B"000000_1000001_00_111",   -- JUMP 65
        
        64 => B"000000000_101_1_01_010", -- MOV R5, AccB
        
        65 => B"000000000_001_0_00_010", -- MOV AccA, R1
        66 => B"000000000_011_0_00_011", -- ADD AccA, R3
        67 => B"000000000_001_0_01_010", -- MOV R1, AccA
        
        68 => B"0_1111001_0_010_0_10_101", -- CNJE R2, AccA, -7
        
        69 => B"000000_1000101_00_111",   -- JUMP 69 (Travado)

        others => B"000000000000000000"
    );
    begin
        dado <= conteudo_rom(to_integer(endereco));
end architecture;